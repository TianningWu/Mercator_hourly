netcdf Mercator_2025-04-25_zos_uovo_6hr {
dimensions:
	time = UNLIMITED ;
	depth = 1 ;
	latitude = 169 ;
	longitude = 289 ;
variables:
	float zos(time, depth, latitude, longitude) ;
		zos:_FillValue = 9.96921e+36f ;
		zos:valid_min = -5.f ;
		zos:valid_max = 5.f ;
		string zos:unit_long = "Meters" ;
		string zos:long_name = "Sea surface height" ;
		string zos:units = "m" ;
		string zos:standard_name = "sea_surface_height_above_geoid" ;
	float uo(time, depth, latitude, longitude) ;
		uo:_FillValue = 9.96921e+36f ;
		uo:valid_min = -10.f ;
		uo:valid_max = 10.f ;
		string uo:unit_long = "Meters per second" ;
		string uo:long_name = "Eastward surface velocity" ;
		string uo:units = "m s-1" ;
		string uo:standard_name = "eastward_sea_water_velocity" ;
	float vo(time, depth, latitude, longitude) ;
		vo:_FillValue = 9.96921e+36f ;
		vo:valid_min = -10.f ;
		vo:valid_max = 10.f ;
		string vo:unit_long = "Meters per second" ;
		string vo:long_name = "Northward surface velocity" ;
		string vo:units = "m s-1" ;
		string vo:standard_name = "northward_sea_water_velocity" ;
	float depth(depth) ;
		string depth:unit_long = "Meters" ;
		string depth:long_name = "Depth" ;
		string depth:units = "m" ;
		string depth:standard_name = "depth" ;
		string depth:positive = "down" ;
		string depth:axis = "Z" ;
	float latitude(latitude) ;
		string latitude:unit_long = "Degrees North" ;
		string latitude:long_name = "Latitude" ;
		string latitude:units = "degrees_north" ;
		string latitude:standard_name = "latitude" ;
		string latitude:axis = "Y" ;
	float longitude(longitude) ;
		string longitude:unit_long = "Degrees East" ;
		string longitude:long_name = "Longitude" ;
		string longitude:units = "degrees_east" ;
		string longitude:standard_name = "longitude" ;
		string longitude:axis = "X" ;
	float time(time) ;
		string time:unit_long = "Hours Since 1950-01-01" ;
		string time:axis = "T" ;
		string time:long_name = "Time" ;
		string time:standard_name = "time" ;
		string time:units = "hours since 1950-01-01" ;
		string time:calendar = "gregorian" ;

// global attributes:
		string :source = "MOI GLO12" ;
		string :credit = "E.U. Copernicus Marine Service Information (CMEMS)" ;
		string :references = "http://marine.copernicus.eu" ;
		string :institution = "Mercator Ocean International" ;
		string :title = "hourly mean fields from Global Ocean Physics Analysis and Forecast updated Daily" ;
		string :producer = "CMEMS - Global Monitoring and Forecasting Centre" ;
		string :Conventions = "CF-1.8" ;
		string :contact = "https://marine.copernicus.eu/contact" ;
		string :copernicusmarine_version = "2.0.1" ;
}
